// ================================================================
// AUTOSA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// AUTOSA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: SA_BLKBOX_SRC0.v
module SA_BLKBOX_SRC0 (
  Y
 );
output Y ;
assign Y = 1'b0;
endmodule
