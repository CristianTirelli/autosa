// ================================================================
// AUTOSA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// AUTOSA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: SA_AUTOSA_RUBIK_fifo.v
`define FORCE_CONTENTION_ASSERTION_RESET_ACTIVE 1'b1
`include "sa_simulate_x_tick.vh"
module SA_AUTOSA_RUBIK_fifo (
      autosa_core_clk
    , autosa_core_rstn
    , idata_prdy
    , idata_pvld
`ifdef FV_RAND_WR_PAUSE
    , idata_pause
`endif
    , idata_pd
    , odata_prdy
    , odata_pvld
    , odata_pd
    , pwrbus_ram_pd
    );
// spyglass disable_block W401 -- clock is not input to module
input autosa_core_clk;
input autosa_core_rstn;
output idata_prdy;
input idata_pvld;
`ifdef FV_RAND_WR_PAUSE
input idata_pause;
`endif
input [255:0] idata_pd;
input odata_prdy;
output odata_pvld;
output [255:0] odata_pd;
input [31:0] pwrbus_ram_pd;
// Master Clock Gating (SLCG)
//
// We gate the clock(s) when idle or stalled.
// This allows us to turn off numerous miscellaneous flops
// that don't get gated during synthesis for one reason or another.
//
// We gate write side and read side separately.
// If the fifo is synchronous, we also gate the ram separately, but if
// -master_clk_gated_unified or -status_reg/-status_logic_reg is specified,
// then we use one clk gate for write, ram, and read.
//
wire autosa_core_clk_mgated_enable; // assigned by code at end of this module
wire autosa_core_clk_mgated; // used only in synchronous fifos
SA_CLK_gate_power autosa_core_clk_mgate( .clk(autosa_core_clk), .reset_(autosa_core_rstn), .clk_en(autosa_core_clk_mgated_enable), .clk_gated(autosa_core_clk_mgated) );
//
// WRITE SIDE
//
// synopsys translate_off
`ifndef SYNTH_LEVEL1_COMPILE
`ifndef SYNTHESIS
wire wr_pause_rand; // random stalling
`endif
`endif
// synopsys translate_on
wire wr_reserving;
reg idata_pvld_in; // registered idata_pvld
reg [255:0] idata_pd_in; // registered idata_pd
reg wr_busy_in; // inputs being held this cycle?
assign idata_prdy = !wr_busy_in;
wire idata_busy_next; // fwd: fifo busy next?
// factor for better timing with distant idata_pvld signal
wire wr_busy_in_next_wr_req_eq_1 = idata_busy_next;
wire wr_busy_in_next_wr_req_eq_0 = (idata_pvld_in && idata_busy_next) && !wr_reserving;
`ifdef FV_RAND_WR_PAUSE
wire wr_busy_in_next = (idata_pvld? wr_busy_in_next_wr_req_eq_1 : wr_busy_in_next_wr_req_eq_0)
                             || idata_pause ;
`else
wire wr_busy_in_next = (idata_pvld? wr_busy_in_next_wr_req_eq_1 : wr_busy_in_next_wr_req_eq_0)
// synopsys translate_off
                            `ifndef SYNTH_LEVEL1_COMPILE
                            `ifndef SYNTHESIS
                            || wr_pause_rand
                            `endif
                            `endif
// synopsys translate_on
                             ;
`endif
wire wr_busy_in_int;
always @( posedge autosa_core_clk or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        idata_pvld_in <= 1'b0;
        wr_busy_in <= 1'b0;
    end else begin
        wr_busy_in <= wr_busy_in_next;
        if ( !wr_busy_in_int ) begin
            idata_pvld_in <= idata_pvld && !wr_busy_in;
        end
//synopsys translate_off
            else if ( wr_busy_in_int ) begin
        end else begin
            idata_pvld_in <= `x_or_0;
        end
//synopsys translate_on
    end
end
always @( posedge autosa_core_clk ) begin
    if ( !wr_busy_in && idata_pvld ) begin
        idata_pd_in <= idata_pd;
    end
//synopsys translate_off
        else if ( !(!wr_busy_in && idata_pvld) ) begin
    end else begin
        idata_pd_in <= {256{`x_or_0}};
    end
//synopsys translate_on
end
reg idata_busy_int; // copy for internal use
assign wr_reserving = idata_pvld_in && !idata_busy_int; // reserving write space?
reg wr_popping; // fwd: write side sees pop?
reg [6:0] idata_count; // write-side count
wire [6:0] wr_count_next_wr_popping = wr_reserving ? idata_count : (idata_count - 1'd1); // spyglass disable W164a W484
wire [6:0] wr_count_next_no_wr_popping = wr_reserving ? (idata_count + 1'd1) : idata_count; // spyglass disable W164a W484
wire [6:0] wr_count_next = wr_popping ? wr_count_next_wr_popping :
                                               wr_count_next_no_wr_popping;
wire wr_count_next_no_wr_popping_is_80 = ( wr_count_next_no_wr_popping == 7'd80 );
wire wr_count_next_is_80 = wr_popping ? 1'b0 :
                                          wr_count_next_no_wr_popping_is_80;
wire [6:0] wr_limit_muxed; // muxed with simulation/emulation overrides
wire [6:0] wr_limit_reg = wr_limit_muxed;
// VCS coverage off
assign idata_busy_next = wr_count_next_is_80 || // busy next cycle?
                          (wr_limit_reg != 7'd0 && // check idata_limit if != 0
                           wr_count_next >= wr_limit_reg) ;
// VCS coverage on
assign wr_busy_in_int = idata_pvld_in && idata_busy_int;
always @( posedge autosa_core_clk_mgated or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        idata_busy_int <= 1'b0;
        idata_count <= 7'd0;
    end else begin
 idata_busy_int <= idata_busy_next;
 if ( wr_reserving ^ wr_popping ) begin
     idata_count <= wr_count_next;
        end
//synopsys translate_off
            else if ( !(wr_reserving ^ wr_popping) ) begin
        end else begin
            idata_count <= {7{`x_or_0}};
        end
//synopsys translate_on
    end
end
wire wr_pushing = wr_reserving; // data pushed same cycle as idata_pvld_in
//
// RAM
//
reg [6:0] idata_adr; // current write address
wire [6:0] odata_adr_p; // read address to use for ram
wire [255:0] odata_pd_p; // read data directly out of ram
wire rd_enable;
wire ore;
wire [31 : 0] pwrbus_ram_pd;
// Adding parameter for fifogen to disable wr/rd contention assertion in ramgen.
// Fifogen handles this by ignoring the data on the ram data out for that cycle.
sa_ram_rwsp_80x256 #(`FORCE_CONTENTION_ASSERTION_RESET_ACTIVE) ram (
      .clk ( autosa_core_clk )
    , .pwrbus_ram_pd ( pwrbus_ram_pd )
    , .wa ( idata_adr )
    , .we ( wr_pushing )
    , .di ( idata_pd_in )
    , .ra ( odata_adr_p )
    , .re ( rd_enable )
    , .dout ( odata_pd_p )
    , .ore ( ore )
    );
// next idata_adr if wr_pushing=1
wire [6:0] wr_adr_next = (idata_adr == 7'd79) ? 7'd0 : (idata_adr + 1'd1); // spyglass disable W484
// spyglass disable_block W484
always @( posedge autosa_core_clk_mgated or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        idata_adr <= 7'd0;
    end else begin
        if ( wr_pushing ) begin
            idata_adr <= wr_adr_next;
        end
//synopsys translate_off
            else if ( !(wr_pushing) ) begin
        end else begin
            idata_adr <= {7{`x_or_0}};
        end
//synopsys translate_on
    end
end
// spyglass enable_block W484
wire rd_popping; // read side doing pop this cycle?
reg [6:0] odata_adr; // current read address
// next read address
wire [6:0] rd_adr_next = (odata_adr == 7'd79) ? 7'd0 : (odata_adr + 1'd1); // spyglass disable W484
assign odata_adr_p = rd_popping ? rd_adr_next : odata_adr; // for ram
// spyglass disable_block W484
always @( posedge autosa_core_clk_mgated or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        odata_adr <= 7'd0;
    end else begin
        if ( rd_popping ) begin
     odata_adr <= rd_adr_next;
        end
//synopsys translate_off
            else if ( !rd_popping ) begin
        end else begin
            odata_adr <= {7{`x_or_0}};
        end
//synopsys translate_on
    end
end
// spyglass enable_block W484
//
// SYNCHRONOUS BOUNDARY
//
always @( posedge autosa_core_clk_mgated or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        wr_popping <= 1'b0;
    end else begin
 wr_popping <= rd_popping;
    end
end
reg rd_pushing;
always @( posedge autosa_core_clk_mgated or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        rd_pushing <= 1'b0;
    end else begin
 rd_pushing <= wr_pushing; // let data go into ram first
    end
end
//
// READ SIDE
//
reg odata_pvld_p; // data out of fifo is valid
reg odata_pvld_int; // internal copy of odata_pvld
assign odata_pvld = odata_pvld_int;
assign rd_popping = odata_pvld_p && !(odata_pvld_int && !odata_prdy);
reg [6:0] odata_count_p; // read-side fifo count
// spyglass disable_block W164a W484
wire [6:0] rd_count_p_next_rd_popping = rd_pushing ? odata_count_p :
                                                                (odata_count_p - 1'd1);
wire [6:0] rd_count_p_next_no_rd_popping = rd_pushing ? (odata_count_p + 1'd1) :
                                                                    odata_count_p;
// spyglass enable_block W164a W484
wire [6:0] rd_count_p_next = rd_popping ? rd_count_p_next_rd_popping :
                                                     rd_count_p_next_no_rd_popping;
wire rd_count_p_next_rd_popping_not_0 = rd_count_p_next_rd_popping != 0;
wire rd_count_p_next_no_rd_popping_not_0 = rd_count_p_next_no_rd_popping != 0;
wire rd_count_p_next_not_0 = rd_popping ? rd_count_p_next_rd_popping_not_0 :
                                              rd_count_p_next_no_rd_popping_not_0;
assign rd_enable = ((rd_count_p_next_not_0) && ((~odata_pvld_p) || rd_popping)); // anytime data's there and not stalled
always @( posedge autosa_core_clk_mgated or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        odata_count_p <= 7'd0;
        odata_pvld_p <= 1'b0;
    end else begin
        if ( rd_pushing || rd_popping ) begin
     odata_count_p <= rd_count_p_next;
        end
//synopsys translate_off
            else if ( !(rd_pushing || rd_popping ) ) begin
        end else begin
            odata_count_p <= {7{`x_or_0}};
        end
//synopsys translate_on
        if ( rd_pushing || rd_popping ) begin
     odata_pvld_p <= (rd_count_p_next_not_0);
        end
//synopsys translate_off
            else if ( !(rd_pushing || rd_popping ) ) begin
        end else begin
            odata_pvld_p <= `x_or_0;
        end
//synopsys translate_on
    end
end
wire rd_req_next = (odata_pvld_p || (odata_pvld_int && !odata_prdy)) ;
always @( posedge autosa_core_clk_mgated or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        odata_pvld_int <= 1'b0;
    end else begin
        odata_pvld_int <= rd_req_next;
    end
end
assign odata_pd = odata_pd_p;
assign ore = rd_popping;
// Master Clock Gating (SLCG) Enables
//
// plusarg for disabling this stuff:
// synopsys translate_off
`ifndef SYNTH_LEVEL1_COMPILE
`ifndef SYNTHESIS
reg master_clk_gating_disabled; initial master_clk_gating_disabled = $test$plusargs( "fifogen_disable_master_clk_gating" ) != 0;
`endif
`endif
// synopsys translate_on
// synopsys translate_off
`ifndef SYNTH_LEVEL1_COMPILE
`ifndef SYNTHESIS
reg wr_pause_rand_dly;
always @( posedge autosa_core_clk or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        wr_pause_rand_dly <= 1'b0;
    end else begin
        wr_pause_rand_dly <= wr_pause_rand;
    end
end
`endif
`endif
// synopsys translate_on
assign autosa_core_clk_mgated_enable = ((wr_reserving || wr_pushing || rd_popping || wr_popping || (idata_pvld_in && !idata_busy_int) || (idata_busy_int != idata_busy_next)) || (rd_pushing || rd_popping || (odata_pvld_int && odata_prdy) || wr_pushing))
                               `ifdef FIFOGEN_MASTER_CLK_GATING_DISABLED
                               || 1'b1
                               `endif
// synopsys translate_off
          `ifndef SYNTH_LEVEL1_COMPILE
          `ifndef SYNTHESIS
                               || master_clk_gating_disabled || (wr_pause_rand != wr_pause_rand_dly)
          `endif
          `endif
// synopsys translate_on
                               ;
// Simulation and Emulation Overrides of wr_limit(s)
//
`ifdef EMU
`ifdef EMU_FIFO_CFG
// Emulation Global Config Override
//
assign wr_limit_muxed = `EMU_FIFO_CFG.SA_AUTOSA_RUBIK_fifo_wr_limit_override ? `EMU_FIFO_CFG.SA_AUTOSA_RUBIK_fifo_wr_limit : 7'd0;
`else
// No Global Override for Emulation
//
assign wr_limit_muxed = 7'd0;
`endif // EMU_FIFO_CFG
`else // !EMU
`ifdef SYNTH_LEVEL1_COMPILE
// No Override for GCS Compiles
//
assign wr_limit_muxed = 7'd0;
`else
`ifdef SYNTHESIS
// No Override for RTL Synthesis
//
assign wr_limit_muxed = 7'd0;
`else
// RTL Simulation Plusarg Override
// VCS coverage off
reg wr_limit_override;
reg [6:0] wr_limit_override_value;
assign wr_limit_muxed = wr_limit_override ? wr_limit_override_value : 7'd0;
`ifdef SA_ARCHPRO
event reinit;
initial begin
    $display("fifogen reinit initial block %m");
    -> reinit;
end
`endif
`ifdef SA_ARCHPRO
always @( reinit ) begin
`else
initial begin
`endif
    wr_limit_override = 0;
    wr_limit_override_value = 0; // to keep viva happy with dangles
    if ( $test$plusargs( "SA_AUTOSA_RUBIK_fifo_wr_limit" ) ) begin
        wr_limit_override = 1;
        $value$plusargs( "SA_AUTOSA_RUBIK_fifo_wr_limit=%d", wr_limit_override_value);
    end
end
// VCS coverage on
`endif
`endif
`endif
// Random Write-Side Stalling
// synopsys translate_off
`ifndef SYNTH_LEVEL1_COMPILE
`ifndef SYNTHESIS
// VCS coverage off
// leda W339 OFF -- Non synthesizable operator
// leda W372 OFF -- Undefined PLI task
// leda W373 OFF -- Undefined PLI function
// leda W599 OFF -- This construct is not supported by Synopsys
// leda W430 OFF -- Initial statement is not synthesizable
// leda W182 OFF -- Illegal statement for synthesis
// leda W639 OFF -- For synthesis, operands of a division or modulo operation need to be constants
// leda DCVER_274_NV OFF -- This system task is not supported by DC
integer stall_probability; // prob of stalling
integer stall_cycles_min; // min cycles to stall
integer stall_cycles_max; // max cycles to stall
integer stall_cycles_left; // stall cycles left
`ifdef SA_ARCHPRO
always @( reinit ) begin
`else
initial begin
`endif
    stall_probability = 0; // no stalling by default
    stall_cycles_min = 1;
    stall_cycles_max = 10;
`ifdef NO_PLI
`else
    if ( $test$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_probability" ) ) begin
        $value$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_probability=%d", stall_probability);
    end else if ( $test$plusargs( "default_fifo_stall_probability" ) ) begin
        $value$plusargs( "default_fifo_stall_probability=%d", stall_probability);
    end
    if ( $test$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_cycles_min" ) ) begin
        $value$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_cycles_min=%d", stall_cycles_min);
    end else if ( $test$plusargs( "default_fifo_stall_cycles_min" ) ) begin
        $value$plusargs( "default_fifo_stall_cycles_min=%d", stall_cycles_min);
    end
    if ( $test$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_cycles_max" ) ) begin
        $value$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_cycles_max=%d", stall_cycles_max);
    end else if ( $test$plusargs( "default_fifo_stall_cycles_max" ) ) begin
        $value$plusargs( "default_fifo_stall_cycles_max=%d", stall_cycles_max);
    end
`endif
    if ( stall_cycles_min < 1 ) begin
        stall_cycles_min = 1;
    end
    if ( stall_cycles_min > stall_cycles_max ) begin
        stall_cycles_max = stall_cycles_min;
    end
end
`ifdef NO_PLI
`else
// randomization globals
`ifdef SIMTOP_RANDOMIZE_STALLS
  always @( `SIMTOP_RANDOMIZE_STALLS.global_stall_event ) begin
    if ( ! $test$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_probability" ) ) stall_probability = `SIMTOP_RANDOMIZE_STALLS.global_stall_fifo_probability;
    if ( ! $test$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_cycles_min" ) ) stall_cycles_min = `SIMTOP_RANDOMIZE_STALLS.global_stall_fifo_cycles_min;
    if ( ! $test$plusargs( "SA_AUTOSA_RUBIK_fifo_fifo_stall_cycles_max" ) ) stall_cycles_max = `SIMTOP_RANDOMIZE_STALLS.global_stall_fifo_cycles_max;
  end
`endif
`endif
always @( negedge autosa_core_clk or negedge autosa_core_rstn ) begin
    if ( !autosa_core_rstn ) begin
        stall_cycles_left <= 0;
    end else begin
`ifdef NO_PLI
            stall_cycles_left <= 0;
`else
            if ( idata_pvld && !(!idata_prdy)
                 && stall_probability != 0 ) begin
                if ( prand_inst0(1, 100) <= stall_probability ) begin
                    stall_cycles_left <= prand_inst1(stall_cycles_min, stall_cycles_max);
                end else if ( stall_cycles_left !== 0 ) begin
                    stall_cycles_left <= stall_cycles_left - 1;
                end
            end else if ( stall_cycles_left !== 0 ) begin
                stall_cycles_left <= stall_cycles_left - 1;
            end
`endif
    end
end
assign wr_pause_rand = (stall_cycles_left !== 0) ;
// VCS coverage on
`endif
`endif
// synopsys translate_on
// VCS coverage on
// leda W339 ON
// leda W372 ON
// leda W373 ON
// leda W599 ON
// leda W430 ON
// leda W182 ON
// leda W639 ON
// leda DCVER_274_NV ON
//
// Histogram of fifo depth (from write side's perspective)
//
// NOTE: it will reference `SIMTOP.perfmon_enabled, so that
// has to at least be defined, though not initialized.
// tbgen testbenches have it already and various
// ways to turn it on and off.
//
`ifdef PERFMON_HISTOGRAM
// synopsys translate_off
`ifndef SYNTH_LEVEL1_COMPILE
`ifndef SYNTHESIS
perfmon_histogram perfmon (
      .clk ( autosa_core_clk )
    , .max ( {25'd0, (wr_limit_reg == 7'd0) ? 7'd80 : wr_limit_reg} )
    , .curr ( {25'd0, idata_count} )
    );
`endif
`endif
// synopsys translate_on
`endif
// spyglass disable_block W164a W164b W116 W484 W504
`ifdef SPYGLASS
`else
`ifdef FV_ASSERT_ON
`else
// synopsys translate_off
`endif
`ifdef ASSERT_ON
`ifdef SPYGLASS
wire disable_assert_plusarg = 1'b0;
`else
`ifdef FV_ASSERT_ON
wire disable_assert_plusarg = 1'b0;
`else
wire disable_assert_plusarg = $test$plusargs("DISABLE_NESS_FLOW_ASSERTIONS");
`endif
`endif
wire assert_enabled = 1'b1 && !disable_assert_plusarg;
`endif
`ifdef FV_ASSERT_ON
`else
// synopsys translate_on
`endif
`ifdef ASSERT_ON
//synopsys translate_off
`ifndef SYNTH_LEVEL1_COMPILE
`ifndef SYNTHESIS
always @(assert_enabled) begin
    if ( assert_enabled === 1'b0 ) begin
        $display("Asserts are disabled for %m");
    end
end
`endif
`endif
//synopsys translate_on
`endif
`endif
// spyglass enable_block W164a W164b W116 W484 W504
//The SA_BLKBOX_SRC0 module is only present when the FIFOGEN_MODULE_SEARCH
// define is set. This is to aid fifogen team search for fifogen fifo
// instance and module names in a given design.
`ifdef FIFOGEN_MODULE_SEARCH
SA_BLKBOX_SRC0 dummy_breadcrumb_fifogen_blkbox (.Y());
`endif
// spyglass enable_block W401 -- clock is not input to module
// synopsys dc_script_begin
// set_boundary_optimization find(design, "SA_AUTOSA_RUBIK_fifo") true
// synopsys dc_script_end
`ifdef SYNTH_LEVEL1_COMPILE
`else
`ifdef SYNTHESIS
`else
`ifdef PRAND_VERILOG
// Only verilog needs any local variables
reg [47:0] prand_local_seed0;
reg prand_initialized0;
reg prand_no_rollpli0;
`endif
`endif
`endif
function [31:0] prand_inst0;
//VCS coverage off
    input [31:0] min;
    input [31:0] max;
    reg [32:0] diff;
    begin
`ifdef SYNTH_LEVEL1_COMPILE
        prand_inst0 = min;
`else
`ifdef SYNTHESIS
        prand_inst0 = min;
`else
`ifdef PRAND_VERILOG
        if (prand_initialized0 !== 1'b1) begin
            prand_no_rollpli0 = $test$plusargs("NO_ROLLPLI");
            if (!prand_no_rollpli0)
                prand_local_seed0 = {$prand_get_seed(0), 16'b0};
            prand_initialized0 = 1'b1;
        end
        if (prand_no_rollpli0) begin
            prand_inst0 = min;
        end else begin
            diff = max - min + 1;
            prand_inst0 = min + prand_local_seed0[47:16] % diff;
// magic numbers taken from Java's random class (same as lrand48)
            prand_local_seed0 = prand_local_seed0 * 48'h5deece66d + 48'd11;
        end
`else
`ifdef PRAND_OFF
        prand_inst0 = min;
`else
        prand_inst0 = $RollPLI(min, max, "auto");
`endif
`endif
`endif
`endif
    end
//VCS coverage on
endfunction
`ifdef SYNTH_LEVEL1_COMPILE
`else
`ifdef SYNTHESIS
`else
`ifdef PRAND_VERILOG
// Only verilog needs any local variables
reg [47:0] prand_local_seed1;
reg prand_initialized1;
reg prand_no_rollpli1;
`endif
`endif
`endif
function [31:0] prand_inst1;
//VCS coverage off
    input [31:0] min;
    input [31:0] max;
    reg [32:0] diff;
    begin
`ifdef SYNTH_LEVEL1_COMPILE
        prand_inst1 = min;
`else
`ifdef SYNTHESIS
        prand_inst1 = min;
`else
`ifdef PRAND_VERILOG
        if (prand_initialized1 !== 1'b1) begin
            prand_no_rollpli1 = $test$plusargs("NO_ROLLPLI");
            if (!prand_no_rollpli1)
                prand_local_seed1 = {$prand_get_seed(1), 16'b0};
            prand_initialized1 = 1'b1;
        end
        if (prand_no_rollpli1) begin
            prand_inst1 = min;
        end else begin
            diff = max - min + 1;
            prand_inst1 = min + prand_local_seed1[47:16] % diff;
// magic numbers taken from Java's random class (same as lrand48)
            prand_local_seed1 = prand_local_seed1 * 48'h5deece66d + 48'd11;
        end
`else
`ifdef PRAND_OFF
        prand_inst1 = min;
`else
        prand_inst1 = $RollPLI(min, max, "auto");
`endif
`endif
`endif
`endif
    end
//VCS coverage on
endfunction
endmodule // SA_AUTOSA_RUBIK_fifo
