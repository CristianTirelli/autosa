// ================================================================
// AUTOSA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// AUTOSA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: SA_AUTOSA_SDP_AUTOSAHLS_X_int_trt.v
module SA_AUTOSA_SDP_AUTOSAHLS_X_int_trt (
   bypass_trt_in //|< i
  ,cfg_mul_shift_value //|< i
  ,mul_data_out //|< i
  ,mul_out_pvld //|< i
  ,autosa_core_clk //|< i
  ,autosa_core_rstn //|< i
  ,trt_out_prdy //|< i
  ,mul_out_prdy //|> o
  ,trt_data_out //|> o
  ,trt_out_pvld //|> o
  );
//parameter X_MUL_OUT_WIDTH = 49;
//parameter X_OUT_WIDTH = 32;
input autosa_core_clk;
input autosa_core_rstn;
input [5:0] cfg_mul_shift_value;
input bypass_trt_in;
input [48:0] mul_data_out;
input mul_out_pvld;
output mul_out_prdy;
output [31:0] trt_data_out;
output trt_out_pvld;
input trt_out_prdy;
reg [31:0] trt_dout;
wire [31:0] trt_data_final;
// synoff nets
// monitor nets
// debug nets
// tie high nets
// tie low nets
// no connect nets
// not all bits used nets
// todo nets
SA_AUTOSA_AUTOSAHLS_shiftrightsu #(.IN_WIDTH(49 ),.OUT_WIDTH(32 ),.SHIFT_WIDTH(6)) x_trt_shiftright_su (
   .data_in ((bypass_trt_in ? 0 : mul_data_out[48:0])) //|< ?
  ,.shift_num (cfg_mul_shift_value[5:0]) //|< i
  ,.data_out (trt_data_final[31:0]) //|> w
  );
//signed
//unsigned
always @(
  bypass_trt_in
  or mul_data_out
  or trt_data_final
  ) begin
   if (bypass_trt_in)
      trt_dout[31:0] = mul_data_out[31:0]; //morework
   else
      trt_dout[31:0] = trt_data_final[31:0];
end
SA_AUTOSA_SDP_AUTOSAHLS_X_INT_TRT_pipe_p1 pipe_p1 (
   .autosa_core_clk (autosa_core_clk) //|< i
  ,.autosa_core_rstn (autosa_core_rstn) //|< i
  ,.mul_out_pvld (mul_out_pvld) //|< i
  ,.trt_dout (trt_dout[31:0]) //|< r
  ,.trt_out_prdy (trt_out_prdy) //|< i
  ,.mul_out_prdy (mul_out_prdy) //|> o
  ,.trt_data_out (trt_data_out[31:0]) //|> o
  ,.trt_out_pvld (trt_out_pvld) //|> o
  );
endmodule // SA_AUTOSA_SDP_AUTOSAHLS_X_int_trt
// **************************************************************************************************************
// Generated by ::pipe -m -bc -rand none -is trt_data_out[31:0] (trt_out_pvld,trt_out_prdy) <= trt_dout[31:0] (mul_out_pvld,mul_out_prdy)
// **************************************************************************************************************
module SA_AUTOSA_SDP_AUTOSAHLS_X_INT_TRT_pipe_p1 (
   autosa_core_clk
  ,autosa_core_rstn
  ,mul_out_pvld
  ,trt_dout
  ,trt_out_prdy
  ,mul_out_prdy
  ,trt_data_out
  ,trt_out_pvld
  );
input autosa_core_clk;
input autosa_core_rstn;
input mul_out_pvld;
input [31:0] trt_dout;
input trt_out_prdy;
output mul_out_prdy;
output [31:0] trt_data_out;
output trt_out_pvld;
reg mul_out_prdy;
reg [31:0] p1_pipe_data;
reg p1_pipe_ready;
reg p1_pipe_ready_bc;
reg p1_pipe_valid;
reg p1_skid_catch;
reg [31:0] p1_skid_data;
reg [31:0] p1_skid_pipe_data;
reg p1_skid_pipe_ready;
reg p1_skid_pipe_valid;
reg p1_skid_ready;
reg p1_skid_ready_flop;
reg p1_skid_valid;
reg [31:0] trt_data_out;
reg trt_out_pvld;
//## pipe (1) skid buffer
always @(
  mul_out_pvld
  or p1_skid_ready_flop
  or p1_skid_pipe_ready
  or p1_skid_valid
  ) begin
  p1_skid_catch = mul_out_pvld && p1_skid_ready_flop && !p1_skid_pipe_ready;
  p1_skid_ready = (p1_skid_valid)? p1_skid_pipe_ready : !p1_skid_catch;
end
always @(posedge autosa_core_clk or negedge autosa_core_rstn) begin
  if (!autosa_core_rstn) begin
    p1_skid_valid <= 1'b0;
    p1_skid_ready_flop <= 1'b1;
    mul_out_prdy <= 1'b1;
  end else begin
  p1_skid_valid <= (p1_skid_valid)? !p1_skid_pipe_ready : p1_skid_catch;
  p1_skid_ready_flop <= p1_skid_ready;
  mul_out_prdy <= p1_skid_ready;
  end
end
always @(posedge autosa_core_clk) begin
// VCS sop_coverage_off start
  p1_skid_data <= (p1_skid_catch)? trt_dout[31:0] : p1_skid_data;
// VCS sop_coverage_off end
end
always @(
  p1_skid_ready_flop
  or mul_out_pvld
  or p1_skid_valid
  or trt_dout
  or p1_skid_data
  ) begin
  p1_skid_pipe_valid = (p1_skid_ready_flop)? mul_out_pvld : p1_skid_valid;
// VCS sop_coverage_off start
  p1_skid_pipe_data = (p1_skid_ready_flop)? trt_dout[31:0] : p1_skid_data;
// VCS sop_coverage_off end
end
//## pipe (1) valid-ready-bubble-collapse
always @(
  p1_pipe_ready
  or p1_pipe_valid
  ) begin
  p1_pipe_ready_bc = p1_pipe_ready || !p1_pipe_valid;
end
always @(posedge autosa_core_clk or negedge autosa_core_rstn) begin
  if (!autosa_core_rstn) begin
    p1_pipe_valid <= 1'b0;
  end else begin
  p1_pipe_valid <= (p1_pipe_ready_bc)? p1_skid_pipe_valid : 1'd1;
  end
end
always @(posedge autosa_core_clk) begin
// VCS sop_coverage_off start
  p1_pipe_data <= (p1_pipe_ready_bc && p1_skid_pipe_valid)? p1_skid_pipe_data : p1_pipe_data;
// VCS sop_coverage_off end
end
always @(
  p1_pipe_ready_bc
  ) begin
  p1_skid_pipe_ready = p1_pipe_ready_bc;
end
//## pipe (1) output
always @(
  p1_pipe_valid
  or trt_out_prdy
  or p1_pipe_data
  ) begin
  trt_out_pvld = p1_pipe_valid;
  p1_pipe_ready = trt_out_prdy;
  trt_data_out[31:0] = p1_pipe_data;
end
//## pipe (1) assertions/testpoints
`ifndef VIVA_PLUGIN_PIPE_DISABLE_ASSERTIONS
wire p1_assert_clk = autosa_core_clk;
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML
// spyglass disable_block STARC-2.10.3.2a
// spyglass disable_block STARC05-2.1.3.1
// spyglass disable_block STARC-2.1.4.6
// spyglass disable_block W116
// spyglass disable_block W154
// spyglass disable_block W239
// spyglass disable_block W362
// spyglass disable_block WRN_58
// spyglass disable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET autosa_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET autosa_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === autosa_core_rstn) ? 1'b0 : autosa_core_rstn)
`else
`define ASSERT_RESET ((1'bx === autosa_core_rstn) ? 1'b1 : autosa_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
`ifndef SYNTHESIS
// VCS coverage off
  sa_assert_no_x #(0,1,0,"No X's allowed on control signals") zzz_assert_no_x_1x (autosa_core_clk, `ASSERT_RESET, autosa_core_rstn, (trt_out_pvld^trt_out_prdy^mul_out_pvld^mul_out_prdy)); // spyglass disable W504 SelfDeterminedExpr-ML 
// VCS coverage on
`endif
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML
// spyglass enable_block STARC-2.10.3.2a
// spyglass enable_block STARC05-2.1.3.1
// spyglass enable_block STARC-2.1.4.6
// spyglass enable_block W116
// spyglass enable_block W154
// spyglass enable_block W239
// spyglass enable_block W362
// spyglass enable_block WRN_58
// spyglass enable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass disable_block NoWidthInBasedNum-ML
// spyglass disable_block STARC-2.10.3.2a
// spyglass disable_block STARC05-2.1.3.1
// spyglass disable_block STARC-2.1.4.6
// spyglass disable_block W116
// spyglass disable_block W154
// spyglass disable_block W239
// spyglass disable_block W362
// spyglass disable_block WRN_58
// spyglass disable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`ifdef ASSERT_ON
`ifdef FV_ASSERT_ON
`define ASSERT_RESET autosa_core_rstn
`else
`ifdef SYNTHESIS
`define ASSERT_RESET autosa_core_rstn
`else
`ifdef ASSERT_OFF_RESET_IS_X
`define ASSERT_RESET ((1'bx === autosa_core_rstn) ? 1'b0 : autosa_core_rstn)
`else
`define ASSERT_RESET ((1'bx === autosa_core_rstn) ? 1'b1 : autosa_core_rstn)
`endif // ASSERT_OFF_RESET_IS_X
`endif // SYNTHESIS
`endif // FV_ASSERT_ON
// VCS coverage off
  sa_assert_hold_throughout_event_interval #(0,1,0,"valid removed before ready") zzz_assert_hold_throughout_event_interval_2x (autosa_core_clk, `ASSERT_RESET, (mul_out_pvld && !mul_out_prdy), (mul_out_pvld), (mul_out_prdy)); // spyglass disable W504 SelfDeterminedExpr-ML 
// VCS coverage on
`undef ASSERT_RESET
`endif // ASSERT_ON
`ifdef SPYGLASS_ASSERT_ON
`else
// spyglass enable_block NoWidthInBasedNum-ML
// spyglass enable_block STARC-2.10.3.2a
// spyglass enable_block STARC05-2.1.3.1
// spyglass enable_block STARC-2.1.4.6
// spyglass enable_block W116
// spyglass enable_block W154
// spyglass enable_block W239
// spyglass enable_block W362
// spyglass enable_block WRN_58
// spyglass enable_block WRN_61
`endif // SPYGLASS_ASSERT_ON
`endif
endmodule // SA_AUTOSA_SDP_AUTOSAHLS_X_INT_TRT_pipe_p1
