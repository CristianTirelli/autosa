// ================================================================
// AUTOSA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// AUTOSA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: SA_AUTOSA_SDP_mrdma.v
// ================================================================
// AUTOSA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// AUTOSA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================
// File Name: SA_AUTOSA_SDP_define.h
module SA_AUTOSA_SDP_mrdma (
   autosa_core_clk //|< i
  ,autosa_core_rstn //|< i
  ,pwrbus_ram_pd //|< i
  ,dla_clk_ovr_on_sync //|< i
  ,global_clk_ovr_on_sync //|< i
  ,tmc2slcg_disable_clock_gating //|< i
  ,mrdma_slcg_op_en //|< i
  ,mrdma_disable //|< i
  ,sdp2mcif_rd_cdt_lat_fifo_pop //|> o
  ,sdp2mcif_rd_req_pd //|> o
  ,sdp2mcif_rd_req_valid //|> o
  ,sdp2mcif_rd_req_ready //|< i
  ,mcif2sdp_rd_rsp_pd //|< i
  ,mcif2sdp_rd_rsp_valid //|< i
  ,mcif2sdp_rd_rsp_ready //|> o
  ,sdp_mrdma2cmux_pd //|> o
  ,sdp_mrdma2cmux_valid //|> o
  ,sdp_mrdma2cmux_ready //|< i
  ,reg2dp_op_en //|< i
  ,reg2dp_batch_number //|< i
  ,reg2dp_channel //|< i
  ,reg2dp_height //|< i
  ,reg2dp_width //|< i
  ,reg2dp_in_precision //|< i
  ,reg2dp_proc_precision //|< i
  ,reg2dp_src_ram_type //|< i
  ,reg2dp_src_base_addr_high //|< i
  ,reg2dp_src_base_addr_low //|< i
  ,reg2dp_src_line_stride //|< i
  ,reg2dp_src_surface_stride //|< i
  ,reg2dp_perf_dma_en //|< i
  ,reg2dp_perf_nan_inf_count_en //|< i
  ,dp2reg_done //|> o
  ,dp2reg_mrdma_stall //|> o
  ,dp2reg_status_inf_input_num //|> o
  ,dp2reg_status_nan_input_num //|> o
  );
//
// SA_AUTOSA_SDP_mrdma_ports.v
//
 input autosa_core_clk;
 input autosa_core_rstn;
 input [31:0] pwrbus_ram_pd;
 input dla_clk_ovr_on_sync;
 input global_clk_ovr_on_sync;
 input tmc2slcg_disable_clock_gating;
 input mrdma_disable;
 input mrdma_slcg_op_en;
 output sdp2mcif_rd_req_valid;
 input sdp2mcif_rd_req_ready;
 output [47 -1:0] sdp2mcif_rd_req_pd;
 input mcif2sdp_rd_rsp_valid;
 output mcif2sdp_rd_rsp_ready;
 input [65 -1:0] mcif2sdp_rd_rsp_pd;
 output sdp2mcif_rd_cdt_lat_fifo_pop;
 output sdp_mrdma2cmux_valid;
 input sdp_mrdma2cmux_ready;
 output [32*8 +1:0] sdp_mrdma2cmux_pd;
 input reg2dp_op_en;
 input [4:0] reg2dp_batch_number;
 input [12:0] reg2dp_channel;
 input [12:0] reg2dp_height;
 input [12:0] reg2dp_width;
 input [1:0] reg2dp_in_precision;
 input [1:0] reg2dp_proc_precision;
 input reg2dp_src_ram_type;
 input [31:0] reg2dp_src_base_addr_high;
 input [31-3:0] reg2dp_src_base_addr_low;
 input [31-3:0] reg2dp_src_line_stride;
 input [31-3:0] reg2dp_src_surface_stride;
 input reg2dp_perf_dma_en;
 input reg2dp_perf_nan_inf_count_en;
 output dp2reg_done;
 output [31:0] dp2reg_mrdma_stall;
 output [31:0] dp2reg_status_inf_input_num;
 output [31:0] dp2reg_status_nan_input_num;
 reg layer_process;
 wire autosa_gated_clk;
 wire op_load;
 wire eg_done;
 wire [13:0] cq2eg_pd;
 wire cq2eg_prdy;
 wire cq2eg_pvld;
 wire [13:0] ig2cq_pd;
 wire ig2cq_prdy;
 wire ig2cq_pvld;
 wire dma_rd_cdt_lat_fifo_pop;
 wire [47 -1:0] dma_rd_req_pd;
 wire dma_rd_req_ram_type;
 wire dma_rd_req_rdy;
 wire dma_rd_req_vld;
 wire dma_rd_rsp_ram_type;
 wire [65 -1:0] dma_rd_rsp_pd;
 wire dma_rd_rsp_rdy;
 wire dma_rd_rsp_vld;
//==============
// Work Processing
//==============
assign op_load = reg2dp_op_en & ~layer_process;
always @(posedge autosa_core_clk or negedge autosa_core_rstn) begin
  if (!autosa_core_rstn) begin
    layer_process <= 1'b0;
  end else begin
    if (op_load) begin
        layer_process <= 1'b1;
    end else if (eg_done) begin
        layer_process <= 1'b0;
    end
  end
end
assign dp2reg_done = eg_done;
//=======================================
 SA_AUTOSA_SDP_MRDMA_gate u_gate (
    .autosa_core_clk (autosa_core_clk) //|< i
   ,.autosa_core_rstn (autosa_core_rstn) //|< i
   ,.dla_clk_ovr_on_sync (dla_clk_ovr_on_sync) //|< i
   ,.global_clk_ovr_on_sync (global_clk_ovr_on_sync) //|< i
   ,.tmc2slcg_disable_clock_gating (tmc2slcg_disable_clock_gating) //|< i
   ,.mrdma_slcg_op_en (mrdma_slcg_op_en) //|< i
   ,.mrdma_disable (mrdma_disable) //|< i
   ,.autosa_gated_clk (autosa_gated_clk) //|> w
   );
//=======================================
// Ingress: send read request to external mem
//---------------------------------------
 SA_AUTOSA_SDP_MRDMA_ig u_ig (
    .autosa_core_clk (autosa_gated_clk) //|< w
   ,.autosa_core_rstn (autosa_core_rstn) //|< i
   ,.op_load (op_load) //|< w
   ,.ig2cq_prdy (ig2cq_prdy) //|< w
   ,.ig2cq_pd (ig2cq_pd[13:0]) //|> w
   ,.ig2cq_pvld (ig2cq_pvld) //|> w
   ,.dma_rd_req_rdy (dma_rd_req_rdy) //|< w
   ,.dma_rd_req_pd (dma_rd_req_pd[47 -1:0]) //|> w
   ,.dma_rd_req_ram_type (dma_rd_req_ram_type) //|> w
   ,.dma_rd_req_vld (dma_rd_req_vld) //|> w
   ,.reg2dp_batch_number (reg2dp_batch_number[4:0]) //|< i
   ,.reg2dp_channel (reg2dp_channel[12:0]) //|< i
   ,.reg2dp_height (reg2dp_height[12:0]) //|< i
   ,.reg2dp_width (reg2dp_width[12:0]) //|< i
   ,.reg2dp_in_precision (reg2dp_in_precision[1:0]) //|< i
   ,.reg2dp_proc_precision (reg2dp_proc_precision[1:0]) //|< i
   ,.reg2dp_src_ram_type (reg2dp_src_ram_type) //|< i
   ,.reg2dp_src_base_addr_high (reg2dp_src_base_addr_high[31:0]) //|< i
   ,.reg2dp_src_base_addr_low (reg2dp_src_base_addr_low[31-3:0]) //|< i
   ,.reg2dp_src_line_stride (reg2dp_src_line_stride[31-3:0]) //|< i
   ,.reg2dp_src_surface_stride (reg2dp_src_surface_stride[31-3:0]) //|< i
   ,.reg2dp_perf_dma_en (reg2dp_perf_dma_en) //|< i
   ,.dp2reg_mrdma_stall (dp2reg_mrdma_stall[31:0]) //|> o
   );
//=======================================
// Context Queue: trace outstanding req, and pass info from Ig to Eg
//---------------------------------------
//: my $depth = (8 < 16) ? 16 : 8;
//: my $width = 14;
//: print "SA_AUTOSA_SDP_MRDMA_cq_${depth}x${width}  u_cq ( \n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
SA_AUTOSA_SDP_MRDMA_cq_16x14  u_cq ( 

//| eperl: generated_end (DO NOT EDIT ABOVE)
    .autosa_core_clk (autosa_gated_clk) //|< w
   ,.autosa_core_rstn (autosa_core_rstn) //|< i
   ,.pwrbus_ram_pd (pwrbus_ram_pd[31:0]) //|< i
   ,.ig2cq_prdy (ig2cq_prdy) //|> w
   ,.ig2cq_pvld (ig2cq_pvld) //|< w
   ,.ig2cq_pd (ig2cq_pd[13:0]) //|< w
   ,.cq2eg_prdy (cq2eg_prdy) //|< w
   ,.cq2eg_pvld (cq2eg_pvld) //|> w
   ,.cq2eg_pd (cq2eg_pd[13:0]) //|> w
   );
//=======================================
// Egress: get return data from external mem
//---------------------------------------
 SA_AUTOSA_SDP_MRDMA_eg u_eg (
    .autosa_core_clk (autosa_gated_clk) //|< w
   ,.autosa_core_rstn (autosa_core_rstn) //|< i
   ,.pwrbus_ram_pd (pwrbus_ram_pd[31:0]) //|< i
   ,.op_load (op_load) //|< w
   ,.eg_done (eg_done) //|> w
   ,.cq2eg_pd (cq2eg_pd[13:0]) //|< w
   ,.cq2eg_pvld (cq2eg_pvld) //|< w
   ,.cq2eg_prdy (cq2eg_prdy) //|> w
   ,.dma_rd_rsp_ram_type (dma_rd_rsp_ram_type) //|> w
   ,.dma_rd_rsp_pd (dma_rd_rsp_pd[65 -1:0]) //|< w
   ,.dma_rd_rsp_rdy (dma_rd_rsp_rdy) //|> w
   ,.dma_rd_rsp_vld (dma_rd_rsp_vld) //|< w
   ,.dma_rd_cdt_lat_fifo_pop (dma_rd_cdt_lat_fifo_pop) //|> w
   ,.sdp_mrdma2cmux_ready (sdp_mrdma2cmux_ready) //|< i
   ,.sdp_mrdma2cmux_pd (sdp_mrdma2cmux_pd[32*8 +1:0]) //|> o
   ,.sdp_mrdma2cmux_valid (sdp_mrdma2cmux_valid) //|> o
   ,.reg2dp_height (reg2dp_height[12:0]) //|< i
   ,.reg2dp_width (reg2dp_width[12:0]) //|< i
   ,.reg2dp_in_precision (reg2dp_in_precision[1:0]) //|< i
   ,.reg2dp_proc_precision (reg2dp_proc_precision[1:0]) //|< i
   ,.reg2dp_src_ram_type (reg2dp_src_ram_type) //|< i
   ,.reg2dp_perf_nan_inf_count_en (reg2dp_perf_nan_inf_count_en) //|< i
   ,.dp2reg_status_inf_input_num (dp2reg_status_inf_input_num[31:0]) //|> o
   ,.dp2reg_status_nan_input_num (dp2reg_status_nan_input_num[31:0]) //|> o
   );
 SA_AUTOSA_SDP_RDMA_dmaif u_SA_AUTOSA_SDP_RDMA_dmaif (
    .autosa_core_clk (autosa_gated_clk) //|< i
   ,.autosa_core_rstn (autosa_core_rstn) //|< i         fixme
   ,.sdp2mcif_rd_cdt_lat_fifo_pop (sdp2mcif_rd_cdt_lat_fifo_pop) //|> o
   ,.sdp2mcif_rd_req_pd (sdp2mcif_rd_req_pd[47 -1:0]) //|> o
   ,.sdp2mcif_rd_req_valid (sdp2mcif_rd_req_valid) //|> o
   ,.sdp2mcif_rd_req_ready (sdp2mcif_rd_req_ready) //|< i
   ,.mcif2sdp_rd_rsp_pd (mcif2sdp_rd_rsp_pd[65 -1:0]) //|< i
   ,.mcif2sdp_rd_rsp_valid (mcif2sdp_rd_rsp_valid) //|< i
   ,.mcif2sdp_rd_rsp_ready (mcif2sdp_rd_rsp_ready) //|> o
   ,.dma_rd_cdt_lat_fifo_pop (dma_rd_cdt_lat_fifo_pop) //|< w
   ,.dma_rd_req_pd (dma_rd_req_pd[47 -1:0]) //|< w
   ,.dma_rd_req_ram_type (dma_rd_req_ram_type) //|< w
   ,.dma_rd_req_vld (dma_rd_req_vld) //|< w
   ,.dma_rd_rsp_ram_type (dma_rd_rsp_ram_type) //|< w
   ,.dma_rd_rsp_rdy (dma_rd_rsp_rdy) //|< w
   ,.dma_rd_req_rdy (dma_rd_req_rdy) //|> w
   ,.dma_rd_rsp_pd (dma_rd_rsp_pd[65 -1:0]) //|> w
   ,.dma_rd_rsp_vld (dma_rd_rsp_vld) //|> w
   );
endmodule // SA_AUTOSA_SDP_mrdma
