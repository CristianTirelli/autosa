// ================================================================
// AUTOSA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// AUTOSA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: SA_BLKBOX_BUFFER.v
module SA_BLKBOX_BUFFER (
  Y
 ,A
 );
output Y ;
input A ;
assign Y = A;
endmodule
